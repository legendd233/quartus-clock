library verilog;
use verilog.vl_types.all;
entity final_vlg_check_tst is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        beep            : in     vl_logic;
        c               : in     vl_logic;
        d               : in     vl_logic;
        e               : in     vl_logic;
        f               : in     vl_logic;
        g               : in     vl_logic;
        h               : in     vl_logic;
        hh              : in     vl_logic;
        j               : in     vl_logic;
        k               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end final_vlg_check_tst;
