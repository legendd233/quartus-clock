library verilog;
use verilog.vl_types.all;
entity final is
    port(
        beep            : out    vl_logic;
        aa              : in     vl_logic;
        a               : out    vl_logic;
        inputb          : in     vl_logic;
        inputa          : in     vl_logic;
        b               : out    vl_logic;
        c               : out    vl_logic;
        d               : out    vl_logic;
        e               : out    vl_logic;
        f               : out    vl_logic;
        g               : out    vl_logic;
        h               : out    vl_logic;
        j               : out    vl_logic;
        k               : out    vl_logic;
        hh              : out    vl_logic
    );
end final;
